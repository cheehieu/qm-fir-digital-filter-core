`timescale 1ns / 100ps

module uart_tb;

   


endmodule // uart_tb
