`timescale 1ns / 100ps

module sasc_brg(/*AUTOARG*/
   // Outputs
   sio_ce, sio_ce_x4,
   // Inputs
   clk, arst_n
   );
   output          sio_ce;      // baud rate
   output          sio_ce_x4;   // baud rate x 4

   input           clk;
   input           arst_n;

   reg             sio_ce;
   reg             sio_ce_x4;
   
   parameter       br_38400_16MHz = 103; // 16e6 / (38400*4) = 104 = 103 + 1
   parameter       br_31250_40MHz = 319; // 40e6 / (31250*4) = 320 = 319 + 1	
   parameter       br_31250_60MHz = 479; // 60e6 / (31250*4) = 480 = 479 + 1
   parameter       br_57600_40MHz = 173; // 40e6 / (57600*4) = 174 = 173 + 1	
   parameter       br_57600_60MHz = 260; // 60e6 / (57600*4) = 261 = 260 + 1	

//`define BRX4pre &{brx4_cntr[6:5],brx4_cntr[2:0]}
//`define BRX4pre &{brx4_cntr[8],brx4_cntr[5:0]}   // 31250 baud rate 40MHz
//`define BRX4pre &{brx4_cntr[7],brx4_cntr[5],brx4_cntr[3:2],brx4_cntr[0]} // 57600 baud rate 40MHz
`define BRX4pre &{brx4_cntr[8],brx4_cntr[2]}   // 57600 baud rate 60MHz

   reg [8:0]       brx4_cntr;
   reg [1:0]       br_cntr;
                   
   always @ (posedge clk or negedge arst_n)
     if (~arst_n)
       brx4_cntr <= 0;
     else if (`BRX4pre)
       brx4_cntr <= 0;
     else
       brx4_cntr <= brx4_cntr + 1'b1;

   always @ (posedge clk or negedge arst_n)
     if (~arst_n)
       br_cntr <= 0;
     else if (`BRX4pre)
       br_cntr <= br_cntr + 1'b1;

   always @ (posedge clk or negedge arst_n)
     if (~arst_n)
       begin
          sio_ce_x4 <= 1'b0;
          sio_ce    <= 1'b0;
       end
     else
       begin
          sio_ce_x4 <= `BRX4pre;
          sio_ce    <= (&br_cntr) & (`BRX4pre);
       end
   
endmodule // sasc_brg
